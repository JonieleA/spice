Title stattement
*M<name> <drain> <gate> <source> <bulk> <model name>
M1 drain gate source 0 2SJ56
.model 2SJ56 PMOS (VTO=1 UO=600 VMAX=2E5 L=2.5u LAMBDA=20m KP=25u)
V1 gate source 5
V2 drain source 5
.DC LIN V2 0 5 .1 V1 LIST 1.5 3
.TEMP 27
.STEP LIN M1 1 3 1 ;$MCE LEVEL;DC Analysis
.PLOT DC ID(M1)
;$SpiceType=AMBIGUOUS
