Title stattement
M1 1 out out 0 $GENERIC_N  
M2 out 2 0 0 $GENERIC_N1
.model $GENERIC_N NMOS(VTO=-2 UO=600 VMAX=2E5 L=2.5u LAMBDA=20m KP=25u W=25u)
.model $GENERIC_N1 NMOS(VTO=1 UO=1000 VMAX=2E5 L=2.5u LAMBDA=20m KP=25u W=25u)
V1 1 0 5
V2 2 0 5
.DC LIN V2 0 5 .01
.TEMP 27
.PLOT DC V(OUT)

;$SpiceType=AMBIGUOUS
