������������� ��� �����
V1 1 0 DC 5
D1 1 0 MyDiod
.MODEL MyDiod D
+(IS=1E-11 N=1 ISR=9E-9 NR=2 RS=0.085 TRS1=0.006 TRS2=1.606E-5 IKF=1 BV=16.825
+TBV1=-5.613E-4 TBV2=-1.687E-7 CJO=1.5E-8 VJ=0.874 M=0.333 EG=1.054 TT=2.303E-7 IBV=3.972E-8)
.OPTIONS GMIN=1E-34
.DC LIN V1 0 2.4 0.01 TEMP LIST -60 25 85
.TEMP 25
.PLOT DC I(D1)
.END

;$SpiceType=AMBIGUOUS
