
V1 1 0 AC 1 0
R1 0 2 4500
C1 2 1 10p
.AC DEC 2500 10K 1E8
.TEMP 27
.PLOT AC VDB(2) VP(2)
;$SpiceType=AMBIGUOUS
