
V1 1 4 SIN (0 15 10k 0 0 30)
D1 0 1 $GENERIC
D2 1 3 $GENERIC
D3 0 4 $GENERIC
D4 4 3 $GENERIC
.model $GENERIC D
R1 3 0 4.5k
C1 3 0 10u

.TRAN 1.5e-007 150U 0 1U 
.TEMP 27
.PLOT TRAN V(R1) V(V1)
;$SpiceType=AMBIGUOUS
