������������ �����������
V1 1 0 SIN(0 3 50 0 0 0)
D1 1 2 MyDiod
R1 2 0 10
.MODEL MyDiod D
+(IS=1E-11 N=1 ISR=9E-9 NR=2 RS=0.085 TRS1=0.006 TRS2=1.606E-5 IKF=1 BV=16.825
+TBV1=-5.613E-4 TBV2=-1.687E-7 CJO=1.5E-8 VJ=0.874 M=0.333 EG=1.054 TT=2.303E-7 IBV=3.972E-8)
.OPTIONS GMIN=1E-34
.TRAN 0.001 50M 0 0.1M 
.TEMP 25
.PLOT TRAN V(R1) V(V1) I(R1)
.END
;$SpiceType=AMBIGUOUS
