
V1 plus 0 10
;$SpiceType=AMBIGUOUS
