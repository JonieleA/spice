
V1 1 0 AC 1 0
R1 2 1 4500
C1 0 2 10p
.AC DEC 250 10K 1E8
.TEMP 27
.PLOT AC VDB(2) VP(2)
;$SpiceType=AMBIGUOUS
