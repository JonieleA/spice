
V1 1 0 PULSE(0 5 0.5u 1n 1n 0.2u 0.5u)
R1 0 2 4500
C1 2 1 10p
.TRAN 6e-008 3U 0 
.TEMP 27
.PLOT TRAN V(1) V(2)
;$SpiceType=AMBIGUOUS
