
R1 1 2 4000
R2 2 0 4000
V1 1 0 DC 9
RL 2 0 8000
.DC LIN V1 0 9 0.1
.TEMP 27
.PLOT DC V(2)
;$SpiceType=AMBIGUOUS
